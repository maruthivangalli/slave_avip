//--------------------------------------------------------------------------------------------
//Module:  Top module
//Description:
//  Consists of Package, run_test;
//--------------------------------------------------------------------------------------------

module top;
  
  //-------------------------------------------------------
  // Importing packages
  //-------------------------------------------------------
  import test_pkg::*;
  import uvm_pkg::*;
  
  //-------------------------------------------------------
  // clock, reset instantiation
  //-------------------------------------------------------
  bit clock;
  bit reset;
  
  //-------------------------------------------------------
  // clock-reset generation
  //-------------------------------------------------------
  always begin
    #10 clock =~ clock;     
  end

  always begin 
    #10 reset=~reset;
  end
  
  //-------------------------------------------------------
  // run_test for simulation
  //-------------------------------------------------------
  initial begin
 //   uvm_config_db #(virtual spi_if)::set(null,"*","vif",in0);
    run_test("base_test");
  end

endmodule

