//--------------------------------------------------------------------------------------------
// Module       : Interface
// Description  : Declaration of pin level signals as logic
//--------------------------------------------------------------------------------------------
interface slave_spi_interface;

  logic sclk;
  logic miso;
  logic mosi;
  logic ss;

endinterface
