//--------------------------------------------------------------------------------------------
// Module       : Slave Driver BFM
// Description  : Connects the slave driver bfm with the driver proxy
//--------------------------------------------------------------------------------------------
module slave_driver_bfm(slave_spi_interface inf);

endmodule
